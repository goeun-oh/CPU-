`timescale 1ns / 1ps

module RV32I_Core (
    input  logic        clk,
    input  logic        reset,
    input  logic [31:0] instrCode,
    output logic        dataWe,
    output logic [31:0] instrMemAddr,
    output logic [31:0] dataAddr,
    output logic [31:0] datawData
);
    logic       regFileWe;
    logic [3:0] aluControl;
    logic aluSrcMuxSel;

    ControlUnit U_ControlUnit (.*);
    DataPath U_DataPath (.*);


endmodule
