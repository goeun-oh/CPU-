`timescale 1ns/1ps

module dataPath(

);
endmodule

module alu(
    input logic [1:0] aluOP,
    input logic [7:0] rd1,
    input logic [7:0] rd2,
    output logic [7:0] 
);
endmodule