`define ADD 4'b0000 // {func7[5], func3}
`define SUB 4'b1000
`define SLL 4'b0001
`define SRL 4'b0101
`define SRA 4'b1101
`define SLT 4'b0010
`define SLTU 4'b0011
`define XOR 4'b0100
`define OR 4'b0110
`define AND 4'b0111

`define OP_TYPE_R 7'b0110011
`define OP_TYPE_L 7'b0000011
`define OP_TYPE_I 7'b0010011
`define OP_TYPE_S 7'b0100011
`define OP_TYPE_B 7'b1100011
`define OP_TYPE_LU 7'b0110111
`define OP_TYPE_AU 7'b0010111 //rd=PC+imm<<12 (12 bit 넘는 주소로 jump 하고 싶을 때 사용)
`define OP_TYPE_J 7'b1101111  //jal, C언어에서 함수호출
`define OP_TYPE_JL 7'b1100111 //jalr, C언어 함수 return 

`define BEQ 3'b000
`define BNE 3'b001
`define BLT 3'b100
`define BGE 3'b101
`define BLTU 3'b110
`define BGEU 3'b111
