module rom(
    input logic [31:0] addr,
    output logic [31:0] rdata
);

    logic [31:0] rom_mem [0:15];

    initial begin
        //rom[x] = 32'b func7_rs2_rs1_f3_rd_opcode; //r-type
        rom_mem[0] = 32'b0000000_00001_00010_000_00100_0110011; //add x4,x2,x1
        rom_mem[1] = 32'b0100000_00001_00010_000_00101_0110011; //sub x5,x2,x1
        rom_mem[2] = 32'b0000000_00001_00010_001_00110_0110011; // sll x6,x2,x1
        rom_mem[3] = 32'b0000000_00001_00010_101_00111_0110011; // srl x7,x2,x1
        rom_mem[4] = 32'b0100000_00001_00010_101_01000_0110011; // sra x8,x2,x1
        rom_mem[5] = 32'b0000000_00001_00010_010_01001_0110011; // slt x9,x2,x1
        rom_mem[6] = 32'b0000000_00001_00010_011_01010_0110011; // sltu x10,x2,x1
        rom_mem[7] = 32'b0000000_00001_00010_100_01011_0110011; // xor x11,x2,x1
        rom_mem[8] = 32'b0000000_00001_00010_110_01100_0110011; // or x12,x2,x1
        rom_mem[9] = 32'b0000000_00001_00010_111_01101_0110011; // and x13,x2,x1
    end

    assign rdata = rom_mem[addr[31:2]]; //4의 배수로 가기위해 하위 2bit 무시
endmodule