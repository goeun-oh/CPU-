`timescale 1ns/1ps

module tb_fndPeriph();



endmodule