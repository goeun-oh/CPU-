module GPI(
    
);

endmodule