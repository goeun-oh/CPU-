`timescale 1ns/1ps

module AXI4_Lite_GPIO(

);

endmodule